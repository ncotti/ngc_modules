class counter_seq_loaded extends counter_sequence_item;
    `uvm_object_utils(counter_seq_loaded)

    function new(string name="");
        super.new();
    endfunction: new
endclass: counter_seq_loaded