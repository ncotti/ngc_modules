class counter_driver extends uvm_component;
    uvm
endclass uvm_component;